-- Copyright (C) 2019  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 19.1.0 Build 670 09/22/2019 SJ Lite Edition
-- Created on Wed Jan 04 09:14:49 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ASM IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Start : IN STD_LOGIC := '0';
        B : IN STD_LOGIC := '0';
        S : OUT STD_LOGIC;
        EDD : OUT STD_LOGIC;
        EDS : OUT STD_LOGIC;
        R : OUT STD_LOGIC;
        CE : OUT STD_LOGIC;
        Clear : OUT STD_LOGIC;
        Rdy : OUT STD_LOGIC
    );
END ASM;	

ARCHITECTURE BEHAVIOR OF ASM IS
    TYPE type_fstate IS (state1,state2,state3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Start,B)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            S <= '0';
            EDD <= '0';
            EDS <= '0';
            R <= '0';
            CE <= '0';
            Clear <= '0';
            Rdy <= '0';
        ELSE
            S <= '0';
            EDD <= '0';
            EDS <= '0';
            R <= '0';
            CE <= '0';
            Clear <= '0';
            Rdy <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF ((Start = '1')) THEN
                        reg_fstate <= state2;
                    ELSIF (NOT((Start = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    EDD <= '1';

                    Clear <= '1';

                    R <= '1';

                    EDS <= '1';
                WHEN state2 =>
                    IF ((B = '1')) THEN
                        reg_fstate <= state3;
                    ELSIF (NOT((B = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    S <= '1';

                    IF (NOT((B = '1'))) THEN
                        EDD <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        EDD <= '0';
                    END IF;

                    Clear <= '1';

                    IF (NOT((B = '1'))) THEN
                        CE <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        CE <= '0';
                    END IF;
                WHEN state3 =>
                    IF ((Start = '1')) THEN
                        reg_fstate <= state3;
                    ELSIF (NOT((Start = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    Rdy <= '1';
                WHEN OTHERS => 
                    S <= 'X';
                    EDD <= 'X';
                    EDS <= 'X';
                    R <= 'X';
                    CE <= 'X';
                    Clear <= 'X';
                    Rdy <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
